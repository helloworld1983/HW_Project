library verilog;
use verilog.vl_types.all;
entity tb_alu32 is
end tb_alu32;
