library verilog;
use verilog.vl_types.all;
entity \_and2\ is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        y               : out    vl_logic
    );
end \_and2\;
