library verilog;
use verilog.vl_types.all;
entity \_inv\ is
    port(
        a               : in     vl_logic;
        y               : out    vl_logic
    );
end \_inv\;
